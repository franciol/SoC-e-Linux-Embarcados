
module niosLab2 (
	clk_clk,
	reset_reset_n,
	stepm_name,
	swx_export);	

	input		clk_clk;
	input		reset_reset_n;
	output	[3:0]	stepm_name;
	input	[3:0]	swx_export;
endmodule
