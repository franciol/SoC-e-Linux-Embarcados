
module niosLab2 (
	clk_clk,
	stepm_export,
	reset_reset_n,
	swx_export);	

	input		clk_clk;
	output	[3:0]	stepm_export;
	input		reset_reset_n;
	input	[3:0]	swx_export;
endmodule
